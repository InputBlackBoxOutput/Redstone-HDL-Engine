module _and(Y, X1, X2);
  input X1, X2;
  output Y;
  
  assign Y = X1&X2;
  
endmodule