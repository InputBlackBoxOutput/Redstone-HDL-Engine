module const(L, H);
    output L, H;

    assign L = 1'b0;
    assign H = 1'b1;
endmodule