module test(input [2:0] A, output [2:0] Y);
    assign Y = &A;
endmodule