module _not(Y, X);
  input X;
  output Y;
  
  assign Y=~X;
endmodule